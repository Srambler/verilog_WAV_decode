library verilog;
use verilog.vl_types.all;
entity reg_config_vlg_tst is
end reg_config_vlg_tst;
